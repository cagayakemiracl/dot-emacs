// Copyright (c) %date% %id% All Rights Reserved.
// $Mail: <%mail%>

module %file-without-ext%(/*AUTOARG*/);
   
endmodule // %file-without-ext%
